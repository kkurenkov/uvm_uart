`ifndef INC_UART_IF
`define INC_UART_IF

interface uart_if ();
  logic         rst;
  logic         tx;
endinterface

`endif